// Module:  bus_arbiter
// Author:  Gheorghe Stefan
// Date:    30.03.2020

module bus_arbiter #(
    parameter PRIORITY_SCHEDULING_ALGORITHM = 0 // Parameter used for selecting between priority scheduling algorithms: 0 for strict priority, 1 for round robin 
)(
    // Server interface

    // Client 1 interface
    
    // Client 2 interface

    // Client 3 interface
    
    // Client 4 interface
);
    
endmodule